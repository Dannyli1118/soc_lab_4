// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0

`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_example
 *
 * This is an example of a (trivially simple) user project,
 * showing how the user project can connect to the logic
 * analyzer, the wishbone bus, and the I/O pads.
 *
 * This project generates an integer count, which is output
 * on the user area GPIO pads (digital output only).  The
 * wishbone connection allows the project to be controlled
 * (start and stop) from the management SoC program.
 *
 * See the testbenches in directory "mprj_counter" for the
 * example programs that drive this user project.  The three
 * testbenches are "io_ports", "la_test1", and "la_test2".
 *
 *-------------------------------------------------------------
 */

module user_proj_example #(
    parameter BITS = 32,
    parameter DELAYS=10
)(
`ifdef USE_POWER_PINS
    inout vccd1,	// User area 1 1.8V supply
    inout vssd1,	// User area 1 digital ground
`endif

    // Wishbone Slave ports (WB MI A)
    input wb_clk_i,
    input wb_rst_i,
    input wbs_stb_i,
    input wbs_cyc_i,
    input wbs_we_i,
    input [3:0] wbs_sel_i,
    input [31:0] wbs_dat_i,
    input [31:0] wbs_adr_i,
    output wbs_ack_o,
    output [31:0] wbs_dat_o,

    // Logic Analyzer Signals
    input  [127:0] la_data_in,
    output [127:0] la_data_out,
    input  [127:0] la_oenb,

    // IOs
    input  [`MPRJ_IO_PADS-1:0] io_in,
    output [`MPRJ_IO_PADS-1:0] io_out,
    output [`MPRJ_IO_PADS-1:0] io_oeb,

    // IRQ
    output [2:0] irq
);
    wire clk;
    wire rst;

    wire [`MPRJ_IO_PADS-1:0] io_in;
    wire [`MPRJ_IO_PADS-1:0] io_out;
    wire [`MPRJ_IO_PADS-1:0] io_oeb;

/////////////////////////////////////////// bram counter read
    wire [3:0] bram_WE0;
    wire bram_EN0;
    //wire [31:0] bram_Di0;
    //wire [31:0] bram_Do0;
    //wire [31:0] bram_A0;
    wire decode;
    wire valid;
    
    reg [3:0] delay_10_counter;
    reg [3:0] next_delay_10_counter; 
    reg [31:0] addr_counter;
    reg [31:0] next_addr_counter;

    assign decode = (wbs_adr_i[31:20] == 12'h380);
    assign valid = decode && wbs_stb_i && wbs_cyc_i;
    assign bram_WE0 = (wbs_we_i && valid) ? 4'b1111 : 4'b0000;
    assign bram_EN0 = 1'b1;
    //assign bram_Di0 = wbs_dat_i;
    assign wbs_ack_o = (delay_10_counter == 4'd10) ? 1'b1 : 1'b0;
    //assign wbs_dat_o = ;

    assign io_out = wbs_dat_o;
    assign io_oeb = !wbs_ack_o;

    always @(posedge wb_clk_i, posedge wb_rst_i) begin
        if (wb_rst_i) begin
            delay_10_counter <= 4'd0;
        end else begin
            delay_10_counter <= next_delay_10_counter;
        end
    end

    always @(*) begin
        if (delay_10_counter == 4'd10) begin
            next_delay_10_counter = 4'd0;
        end else if (valid && wbs_ack_o == 1'b0) begin
            next_delay_10_counter = delay_10_counter + 4'd1;
        end else begin
            next_delay_10_counter = delay_10_counter;
        end
    end

    bram user_bram (
        .CLK(wb_clk_i),
        .WE0(bram_WE0),
        .EN0(bram_EN0),
        .Di0(wbs_dat_i),
        .Do0(wbs_dat_o),
        .A0(wbs_adr_i)
    );

endmodule



`default_nettype wire
